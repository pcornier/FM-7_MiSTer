
module m139(
  input clk,
  input [8:0] addr,
  output reg [3:0] q,
  input cs_n,
  output rdy_n
);

  reg old_cs;
  assign rdy_n = old_cs != cs_n;

  always @(posedge clk) begin
    old_cs <= cs_n;
    if (~cs_n) begin
      case (addr)
        9'h000 : q <= 4'h7;
        9'h001 : q <= 4'h7;
        9'h002 : q <= 4'h7;
        9'h003 : q <= 4'h7;
        9'h004 : q <= 4'h7;
        9'h005 : q <= 4'h7;
        9'h006 : q <= 4'h7;
        9'h007 : q <= 4'h7;
        9'h008 : q <= 4'h7;
        9'h009 : q <= 4'h7;
        9'h00a : q <= 4'h7;
        9'h00b : q <= 4'h7;
        9'h00c : q <= 4'h7;
        9'h00d : q <= 4'h7;
        9'h00e : q <= 4'h7;
        9'h00f : q <= 4'h7;
        9'h010 : q <= 4'h7;
        9'h011 : q <= 4'h7;
        9'h012 : q <= 4'h7;
        9'h013 : q <= 4'h7;
        9'h014 : q <= 4'h7;
        9'h015 : q <= 4'h7;
        9'h016 : q <= 4'h7;
        9'h017 : q <= 4'h7;
        9'h018 : q <= 4'h7;
        9'h019 : q <= 4'h7;
        9'h01a : q <= 4'h7;
        9'h01b : q <= 4'h7;
        9'h01c : q <= 4'h7;
        9'h01d : q <= 4'h7;
        9'h01e : q <= 4'h7;
        9'h01f : q <= 4'h7;
        9'h020 : q <= 4'h7;
        9'h021 : q <= 4'h7;
        9'h022 : q <= 4'h7;
        9'h023 : q <= 4'h7;
        9'h024 : q <= 4'h7;
        9'h025 : q <= 4'h7;
        9'h026 : q <= 4'h7;
        9'h027 : q <= 4'h7;
        9'h028 : q <= 4'h7;
        9'h029 : q <= 4'h7;
        9'h02a : q <= 4'h7;
        9'h02b : q <= 4'h7;
        9'h02c : q <= 4'h7;
        9'h02d : q <= 4'h7;
        9'h02e : q <= 4'h7;
        9'h02f : q <= 4'h7;
        9'h030 : q <= 4'h7;
        9'h031 : q <= 4'h7;
        9'h032 : q <= 4'h7;
        9'h033 : q <= 4'h7;
        9'h034 : q <= 4'h7;
        9'h035 : q <= 4'h7;
        9'h036 : q <= 4'h7;
        9'h037 : q <= 4'h7;
        9'h038 : q <= 4'h7;
        9'h039 : q <= 4'h7;
        9'h03a : q <= 4'h7;
        9'h03b : q <= 4'h7;
        9'h03c : q <= 4'h7;
        9'h03d : q <= 4'h7;
        9'h03e : q <= 4'h7;
        9'h03f : q <= 4'h7;
        9'h040 : q <= 4'he;
        9'h041 : q <= 4'he;
        9'h042 : q <= 4'he;
        9'h043 : q <= 4'he;
        9'h044 : q <= 4'he;
        9'h045 : q <= 4'he;
        9'h046 : q <= 4'he;
        9'h047 : q <= 4'he;
        9'h048 : q <= 4'he;
        9'h049 : q <= 4'he;
        9'h04a : q <= 4'he;
        9'h04b : q <= 4'he;
        9'h04c : q <= 4'he;
        9'h04d : q <= 4'he;
        9'h04e : q <= 4'he;
        9'h04f : q <= 4'he;
        9'h050 : q <= 4'he;
        9'h051 : q <= 4'he;
        9'h052 : q <= 4'he;
        9'h053 : q <= 4'he;
        9'h054 : q <= 4'he;
        9'h055 : q <= 4'he;
        9'h056 : q <= 4'he;
        9'h057 : q <= 4'he;
        9'h058 : q <= 4'he;
        9'h059 : q <= 4'he;
        9'h05a : q <= 4'he;
        9'h05b : q <= 4'he;
        9'h05c : q <= 4'he;
        9'h05d : q <= 4'he;
        9'h05e : q <= 4'he;
        9'h05f : q <= 4'he;
        9'h060 : q <= 4'he;
        9'h061 : q <= 4'he;
        9'h062 : q <= 4'he;
        9'h063 : q <= 4'he;
        9'h064 : q <= 4'he;
        9'h065 : q <= 4'he;
        9'h066 : q <= 4'he;
        9'h067 : q <= 4'he;
        9'h068 : q <= 4'he;
        9'h069 : q <= 4'he;
        9'h06a : q <= 4'he;
        9'h06b : q <= 4'he;
        9'h06c : q <= 4'he;
        9'h06d : q <= 4'he;
        9'h06e : q <= 4'he;
        9'h06f : q <= 4'he;
        9'h070 : q <= 4'he;
        9'h071 : q <= 4'he;
        9'h072 : q <= 4'he;
        9'h073 : q <= 4'he;
        9'h074 : q <= 4'he;
        9'h075 : q <= 4'he;
        9'h076 : q <= 4'he;
        9'h077 : q <= 4'he;
        9'h078 : q <= 4'he;
        9'h079 : q <= 4'he;
        9'h07a : q <= 4'he;
        9'h07b : q <= 4'he;
        9'h07c : q <= 4'he;
        9'h07d : q <= 4'he;
        9'h07e : q <= 4'he;
        9'h07f : q <= 4'he;
        9'h080 : q <= 4'hd; // f
        9'h081 : q <= 4'hd; // f
        9'h082 : q <= 4'hd; // f
        9'h083 : q <= 4'hd;
        9'h084 : q <= 4'hd;
        9'h085 : q <= 4'hd;
        9'h086 : q <= 4'hd;
        9'h087 : q <= 4'hd; // f
        9'h088 : q <= 4'hd;
        9'h089 : q <= 4'hd;
        9'h08a : q <= 4'hd;
        9'h08b : q <= 4'hd;
        9'h08c : q <= 4'hd;
        9'h08d : q <= 4'hd;
        9'h08e : q <= 4'hd;
        9'h08f : q <= 4'hd;
        9'h090 : q <= 4'hd;
        9'h091 : q <= 4'hd;
        9'h092 : q <= 4'hd;
        9'h093 : q <= 4'hd;
        9'h094 : q <= 4'hd;
        9'h095 : q <= 4'hd;
        9'h096 : q <= 4'hd; // f
        9'h097 : q <= 4'hd; // f
        9'h098 : q <= 4'hd;
        9'h099 : q <= 4'hd;
        9'h09a : q <= 4'hd;
        9'h09b : q <= 4'hd; // f
        9'h09c : q <= 4'hd; // f
        9'h09d : q <= 4'hd; // f
        9'h09e : q <= 4'hd; // f
        9'h09f : q <= 4'hd; // f
        9'h0a0 : q <= 4'hd;
        9'h0a1 : q <= 4'hd;
        9'h0a2 : q <= 4'hd;
        9'h0a3 : q <= 4'hd;
        9'h0a4 : q <= 4'hd;
        9'h0a5 : q <= 4'hd;
        9'h0a6 : q <= 4'hd;
        9'h0a7 : q <= 4'hd;
        9'h0a8 : q <= 4'hd;
        9'h0a9 : q <= 4'hd;
        9'h0aa : q <= 4'hd;
        9'h0ab : q <= 4'hd;
        9'h0ac : q <= 4'hd;
        9'h0ad : q <= 4'hd;
        9'h0ae : q <= 4'hd;
        9'h0af : q <= 4'hd;
        9'h0b0 : q <= 4'hd;
        9'h0b1 : q <= 4'hd;
        9'h0b2 : q <= 4'hd;
        9'h0b3 : q <= 4'hd;
        9'h0b4 : q <= 4'hd;
        9'h0b5 : q <= 4'hd;
        9'h0b6 : q <= 4'hd;
        9'h0b7 : q <= 4'hd;
        9'h0b8 : q <= 4'hd;
        9'h0b9 : q <= 4'hd;
        9'h0ba : q <= 4'hd;
        9'h0bb : q <= 4'hd;
        9'h0bc : q <= 4'hd;
        9'h0bd : q <= 4'hd;
        9'h0be : q <= 4'hd;
        9'h0bf : q <= 4'hd;
        9'h0c0 : q <= 4'hd;
        9'h0c1 : q <= 4'hd;
        9'h0c2 : q <= 4'hd;
        9'h0c3 : q <= 4'hd;
        9'h0c4 : q <= 4'hd;
        9'h0c5 : q <= 4'hd;
        9'h0c6 : q <= 4'hd;
        9'h0c7 : q <= 4'hd;
        9'h0c8 : q <= 4'hd;
        9'h0c9 : q <= 4'hd;
        9'h0ca : q <= 4'hd;
        9'h0cb : q <= 4'hd;
        9'h0cc : q <= 4'hd;
        9'h0cd : q <= 4'hd;
        9'h0ce : q <= 4'hd;
        9'h0cf : q <= 4'hd;
        9'h0d0 : q <= 4'hd;
        9'h0d1 : q <= 4'hd;
        9'h0d2 : q <= 4'hd;
        9'h0d3 : q <= 4'hd;
        9'h0d4 : q <= 4'hd;
        9'h0d5 : q <= 4'hd;
        9'h0d6 : q <= 4'hd;
        9'h0d7 : q <= 4'hd;
        9'h0d8 : q <= 4'hd;
        9'h0d9 : q <= 4'hd;
        9'h0da : q <= 4'hd;
        9'h0db : q <= 4'hd;
        9'h0dc : q <= 4'hd;
        9'h0dd : q <= 4'hd;
        9'h0de : q <= 4'hd;
        9'h0df : q <= 4'hd;
        9'h0e0 : q <= 4'hd;
        9'h0e1 : q <= 4'hd;
        9'h0e2 : q <= 4'hd;
        9'h0e3 : q <= 4'hd;
        9'h0e4 : q <= 4'hd;
        9'h0e5 : q <= 4'hd;
        9'h0e6 : q <= 4'hd;
        9'h0e7 : q <= 4'hd;
        9'h0e8 : q <= 4'hd;
        9'h0e9 : q <= 4'hd;
        9'h0ea : q <= 4'hd;
        9'h0eb : q <= 4'hd;
        9'h0ec : q <= 4'hd;
        9'h0ed : q <= 4'hd;
        9'h0ee : q <= 4'hd;
        9'h0ef : q <= 4'hd;
        9'h0f0 : q <= 4'hd;
        9'h0f1 : q <= 4'hd;
        9'h0f2 : q <= 4'hd;
        9'h0f3 : q <= 4'hd;
        9'h0f4 : q <= 4'hd;
        9'h0f5 : q <= 4'hd;
        9'h0f6 : q <= 4'hd;
        9'h0f7 : q <= 4'hd;
        9'h0f8 : q <= 4'hd;
        9'h0f9 : q <= 4'hd;
        9'h0fa : q <= 4'hd;
        9'h0fb : q <= 4'hd;
        9'h0fc : q <= 4'hd;
        9'h0fd : q <= 4'hd;
        9'h0fe : q <= 4'hd;
        9'h0ff : q <= 4'hd;
        9'h100 : q <= 4'hb;
        9'h101 : q <= 4'hb;
        9'h102 : q <= 4'hb;
        9'h103 : q <= 4'hb;
        9'h104 : q <= 4'hb;
        9'h105 : q <= 4'hb;
        9'h106 : q <= 4'hb;
        9'h107 : q <= 4'hb;
        9'h108 : q <= 4'hb;
        9'h109 : q <= 4'hb;
        9'h10a : q <= 4'hb;
        9'h10b : q <= 4'hb;
        9'h10c : q <= 4'hb;
        9'h10d : q <= 4'hb;
        9'h10e : q <= 4'hb;
        9'h10f : q <= 4'hb;
        9'h110 : q <= 4'hb;
        9'h111 : q <= 4'hb;
        9'h112 : q <= 4'hb;
        9'h113 : q <= 4'hb;
        9'h114 : q <= 4'hb;
        9'h115 : q <= 4'hb;
        9'h116 : q <= 4'hb;
        9'h117 : q <= 4'hb;
        9'h118 : q <= 4'hb;
        9'h119 : q <= 4'hb;
        9'h11a : q <= 4'hb;
        9'h11b : q <= 4'hb;
        9'h11c : q <= 4'hb;
        9'h11d : q <= 4'hb;
        9'h11e : q <= 4'hb;
        9'h11f : q <= 4'hb;
        9'h120 : q <= 4'hb;
        9'h121 : q <= 4'hb;
        9'h122 : q <= 4'hb;
        9'h123 : q <= 4'hb;
        9'h124 : q <= 4'hb;
        9'h125 : q <= 4'hb;
        9'h126 : q <= 4'hb;
        9'h127 : q <= 4'hb;
        9'h128 : q <= 4'hb;
        9'h129 : q <= 4'hb;
        9'h12a : q <= 4'hb;
        9'h12b : q <= 4'hb;
        9'h12c : q <= 4'hb;
        9'h12d : q <= 4'hb;
        9'h12e : q <= 4'hb;
        9'h12f : q <= 4'hb;
        9'h130 : q <= 4'hb;
        9'h131 : q <= 4'hb;
        9'h132 : q <= 4'hb;
        9'h133 : q <= 4'hb;
        9'h134 : q <= 4'hb;
        9'h135 : q <= 4'hb;
        9'h136 : q <= 4'hb;
        9'h137 : q <= 4'hb;
        9'h138 : q <= 4'hb;
        9'h139 : q <= 4'hb;
        9'h13a : q <= 4'hb;
        9'h13b : q <= 4'hb;
        9'h13c : q <= 4'hb;
        9'h13d : q <= 4'hb;
        9'h13e : q <= 4'hb;
        9'h13f : q <= 4'hb;
        9'h140 : q <= 4'hb;
        9'h141 : q <= 4'hb;
        9'h142 : q <= 4'hb;
        9'h143 : q <= 4'hb;
        9'h144 : q <= 4'hb;
        9'h145 : q <= 4'hb;
        9'h146 : q <= 4'hb;
        9'h147 : q <= 4'hb;
        9'h148 : q <= 4'hb;
        9'h149 : q <= 4'hb;
        9'h14a : q <= 4'hb;
        9'h14b : q <= 4'hb;
        9'h14c : q <= 4'hb;
        9'h14d : q <= 4'hb;
        9'h14e : q <= 4'hb;
        9'h14f : q <= 4'hb;
        9'h150 : q <= 4'hb;
        9'h151 : q <= 4'hb;
        9'h152 : q <= 4'hb;
        9'h153 : q <= 4'hb;
        9'h154 : q <= 4'hb;
        9'h155 : q <= 4'hb;
        9'h156 : q <= 4'hb;
        9'h157 : q <= 4'hb;
        9'h158 : q <= 4'hb;
        9'h159 : q <= 4'hb;
        9'h15a : q <= 4'hb;
        9'h15b : q <= 4'hb;
        9'h15c : q <= 4'hb;
        9'h15d : q <= 4'hb;
        9'h15e : q <= 4'hb;
        9'h15f : q <= 4'hb;
        9'h160 : q <= 4'hb;
        9'h161 : q <= 4'hb;
        9'h162 : q <= 4'hb;
        9'h163 : q <= 4'hb;
        9'h164 : q <= 4'hb;
        9'h165 : q <= 4'hb;
        9'h166 : q <= 4'hb;
        9'h167 : q <= 4'hb;
        9'h168 : q <= 4'hb;
        9'h169 : q <= 4'hb;
        9'h16a : q <= 4'hb;
        9'h16b : q <= 4'hb;
        9'h16c : q <= 4'hb;
        9'h16d : q <= 4'hb;
        9'h16e : q <= 4'hb;
        9'h16f : q <= 4'hb;
        9'h170 : q <= 4'hb;
        9'h171 : q <= 4'hb;
        9'h172 : q <= 4'hb;
        9'h173 : q <= 4'hb;
        9'h174 : q <= 4'hb;
        9'h175 : q <= 4'hb;
        9'h176 : q <= 4'hb;
        9'h177 : q <= 4'hb;
        9'h178 : q <= 4'hb;
        9'h179 : q <= 4'hb;
        9'h17a : q <= 4'hb;
        9'h17b : q <= 4'hb;
        9'h17c : q <= 4'hb;
        9'h17d : q <= 4'hb;
        9'h17e : q <= 4'hb;
        9'h17f : q <= 4'hb;
        9'h180 : q <= 4'hb;
        9'h181 : q <= 4'hb;
        9'h182 : q <= 4'hb;
        9'h183 : q <= 4'hb;
        9'h184 : q <= 4'hb;
        9'h185 : q <= 4'hb;
        9'h186 : q <= 4'hb;
        9'h187 : q <= 4'hb;
        9'h188 : q <= 4'hb;
        9'h189 : q <= 4'hb;
        9'h18a : q <= 4'hb;
        9'h18b : q <= 4'hb;
        9'h18c : q <= 4'hb;
        9'h18d : q <= 4'hb;
        9'h18e : q <= 4'hb;
        9'h18f : q <= 4'hb;
        9'h190 : q <= 4'hb;
        9'h191 : q <= 4'hb;
        9'h192 : q <= 4'hb;
        9'h193 : q <= 4'hb;
        9'h194 : q <= 4'hb;
        9'h195 : q <= 4'hb;
        9'h196 : q <= 4'hb;
        9'h197 : q <= 4'hb;
        9'h198 : q <= 4'hb;
        9'h199 : q <= 4'hb;
        9'h19a : q <= 4'hb;
        9'h19b : q <= 4'hb;
        9'h19c : q <= 4'hb;
        9'h19d : q <= 4'hb;
        9'h19e : q <= 4'hb;
        9'h19f : q <= 4'hb;
        9'h1a0 : q <= 4'hb;
        9'h1a1 : q <= 4'hb;
        9'h1a2 : q <= 4'hb;
        9'h1a3 : q <= 4'hb;
        9'h1a4 : q <= 4'hb;
        9'h1a5 : q <= 4'hb;
        9'h1a6 : q <= 4'hb;
        9'h1a7 : q <= 4'hb;
        9'h1a8 : q <= 4'hb;
        9'h1a9 : q <= 4'hb;
        9'h1aa : q <= 4'hb;
        9'h1ab : q <= 4'hb;
        9'h1ac : q <= 4'hb;
        9'h1ad : q <= 4'hb;
        9'h1ae : q <= 4'hb;
        9'h1af : q <= 4'hb;
        9'h1b0 : q <= 4'hb;
        9'h1b1 : q <= 4'hb;
        9'h1b2 : q <= 4'hb;
        9'h1b3 : q <= 4'hb;
        9'h1b4 : q <= 4'hb;
        9'h1b5 : q <= 4'hb;
        9'h1b6 : q <= 4'hb;
        9'h1b7 : q <= 4'hb;
        9'h1b8 : q <= 4'hb;
        9'h1b9 : q <= 4'hb;
        9'h1ba : q <= 4'hb;
        9'h1bb : q <= 4'hb;
        9'h1bc : q <= 4'hb;
        9'h1bd : q <= 4'hb;
        9'h1be : q <= 4'hb;
        9'h1bf : q <= 4'hb;
        9'h1c0 : q <= 4'hb;
        9'h1c1 : q <= 4'hb;
        9'h1c2 : q <= 4'hb;
        9'h1c3 : q <= 4'hb;
        9'h1c4 : q <= 4'hb;
        9'h1c5 : q <= 4'hb;
        9'h1c6 : q <= 4'hb;
        9'h1c7 : q <= 4'hb;
        9'h1c8 : q <= 4'hb;
        9'h1c9 : q <= 4'hb;
        9'h1ca : q <= 4'hb;
        9'h1cb : q <= 4'hb;
        9'h1cc : q <= 4'hb;
        9'h1cd : q <= 4'hb;
        9'h1ce : q <= 4'hb;
        9'h1cf : q <= 4'hb;
        9'h1d0 : q <= 4'hb;
        9'h1d1 : q <= 4'hb;
        9'h1d2 : q <= 4'hb;
        9'h1d3 : q <= 4'hb;
        9'h1d4 : q <= 4'hb;
        9'h1d5 : q <= 4'hb;
        9'h1d6 : q <= 4'hb;
        9'h1d7 : q <= 4'hb;
        9'h1d8 : q <= 4'hb;
        9'h1d9 : q <= 4'hb;
        9'h1da : q <= 4'hb;
        9'h1db : q <= 4'hb;
        9'h1dc : q <= 4'hb;
        9'h1dd : q <= 4'hb;
        9'h1de : q <= 4'hb;
        9'h1df : q <= 4'hb;
        9'h1e0 : q <= 4'hb;
        9'h1e1 : q <= 4'hb;
        9'h1e2 : q <= 4'hb;
        9'h1e3 : q <= 4'hb;
        9'h1e4 : q <= 4'hb;
        9'h1e5 : q <= 4'hb;
        9'h1e6 : q <= 4'hb;
        9'h1e7 : q <= 4'hb;
        9'h1e8 : q <= 4'hb;
        9'h1e9 : q <= 4'hb;
        9'h1ea : q <= 4'hb;
        9'h1eb : q <= 4'hb;
        9'h1ec : q <= 4'hb;
        9'h1ed : q <= 4'hb;
        9'h1ee : q <= 4'hb;
        9'h1ef : q <= 4'hb;
        9'h1f0 : q <= 4'h7;
        9'h1f1 : q <= 4'h7;
        9'h1f2 : q <= 4'h7;
        9'h1f3 : q <= 4'h7;
        9'h1f4 : q <= 4'h7;
        9'h1f5 : q <= 4'h7;
        9'h1f6 : q <= 4'h7;
        9'h1f7 : q <= 4'h7;
        9'h1f8 : q <= 4'h7;
        9'h1f9 : q <= 4'h7;
        9'h1fa : q <= 4'h7;
        9'h1fb : q <= 4'h7;
        9'h1fc : q <= 4'h7;
        9'h1fd : q <= 4'h7;
        9'h1fe : q <= 4'hb;
        9'h1ff : q <= 4'hb;
        default: q <= 4'h0;
      endcase
    end
    else begin
      q <= 4'h0;
    end
  end

endmodule
